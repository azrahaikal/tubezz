library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;


entity counter is
	port(	clk, rst: in std_logic;
			rstCounter : in std_logic;
			enCounter : in std_logic;
			counterOut : out std_logic_vector(3 downto 0);
			counterOut2 : in std_logic_vector(3 downto 0)
	);
end entity;

architecture counter_arc of counter is
begin
	process(rst, clk, enCounter, counterOut2)
	begin
	if (rst = '1' or rstCounter = '1') then
		counterOut <= "1101";
	elsif (clk'EVENT and clk = '1') then
		if (enCounter = '1') then 
	
		if (counterOut2 = "0000") then
			counterOut <= "0001";
		elsif (counterOut2 = "0001") then
			counterOut <= "0010";
		elsif (counterOut2 = "0010") then
			counterOut <= "0011";
		elsif (counterOut2 = "0011") then
			counterOut <= "0100";
		elsif (counterOut2 = "0100") then
			counterOut <= "0101";
		elsif (counterOut2 = "0101") then
			counterOut <= "0110";
		elsif (counterOut2 = "0110") then
			counterOut <= "0111";
		elsif (counterOut2 = "0111") then
			counterOut <= "1000";
		elsif (counterOut2 = "1000") then
			counterOut <= "1001";
		elsif (counterOut2 = "1001") then
			counterOut <= "1010";
		elsif (counterOut2 = "1010") then
			counterOut <= "1011";
		elsif (counterOut2 = "1011") then
			counterOut <= "1100";
		elsif (counterOut2 = "1100") then
			counterOut <= "1101";
		elsif (counterOut2 = "1101") then
			counterOut <= "0000";
		else
			counterOut <= "1101";			
		end if;
		end if;
	end if;
	end process;
end counter_arc;